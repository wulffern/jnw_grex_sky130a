*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/JNW_GREX_lpe.spi
#else
.include ../../../work/xsch/JNW_GREX.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  VSS  pwl 0 0 10n {AVDD}
VPWR  PWRUP_1V8  VSS  pwl 0 0 1u 0 1.01u {AVDD}
VRESET  RESET_1V8  VSS  pwl 0 {AVDD} 2u {AVDD} 2.01u 0

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save v(do_1v8)
.save v(pwrup_1v8)
.save v(reset_1v8)
.save v(pulse_1v8) v(vdd_1v8) i(vdd) i(vss)
.save v(xdut.iptn) v(xdut.XA_TI1.IPTN) v(xdut.vo_1v8) v(xdut.xa_ti.vbn1) v(xdut.xa_ti.vbn2)
.save all


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0


set fend = .raw
foreach vtemp -40 -20 0 20 40 60 80 100
  option temp=$vtemp
  tran 10n 5u
  write {cicname}_$vtemp$fend
end
quit


.endc

.end
