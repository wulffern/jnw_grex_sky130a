magic
tech sky130A
magscale 1 2
timestamp 1735577829
<< locali >>
rect -3500 6600 2100 7000
rect -3500 1100 -3100 6600
rect -2912 1100 -2720 2196
rect -1888 1100 -1696 2196
rect -1312 1600 -1120 2180
rect -288 1600 -96 2196
rect 388 1600 580 2196
rect 1412 1600 1604 2196
rect -1312 1490 1700 1600
rect -1312 1482 -922 1490
rect -1580 1476 -922 1482
rect -1580 1325 -1575 1476
rect -1424 1325 -922 1476
rect -1580 1319 -922 1325
rect -1312 1310 -922 1319
rect -742 1310 778 1490
rect 958 1393 1700 1490
rect 958 1310 1055 1393
rect -1312 1305 1055 1310
rect 1143 1305 1700 1393
rect -1312 1204 1700 1305
rect -1300 1200 1700 1204
rect 1800 1100 2100 6600
rect -3500 1090 2100 1100
rect -3500 910 -2522 1090
rect -2342 910 2100 1090
rect -3500 900 2100 910
<< viali >>
rect -2475 5924 -2324 6075
rect 1010 6010 1190 6190
rect -1575 1325 -1424 1476
rect -922 1310 -742 1490
rect 778 1310 958 1490
rect 1055 1305 1143 1393
rect -2522 910 -2342 1090
<< metal1 >>
rect 1004 6190 1196 6202
rect -2481 6081 -2318 6087
rect -2481 5912 -2318 5918
rect -1581 6081 -1418 6087
rect -2272 4996 -2080 5002
rect -2656 2932 -2592 2938
rect -2656 2668 -2592 2868
rect -2272 2596 -2080 4804
rect -2528 1090 -2336 2396
rect -1581 1476 -1418 5918
rect 1004 6010 1010 6190
rect 1190 6010 1196 6190
rect 1004 5500 1196 6010
rect 1000 5300 2100 5500
rect 1004 5012 1196 5300
rect 990 4996 1227 5012
rect 990 4804 1004 4996
rect 1196 4804 1227 4996
rect 990 4791 1227 4804
rect 1900 4300 2098 4400
rect 1800 4285 2098 4300
rect 1800 4114 1914 4285
rect 2085 4114 2098 4285
rect 1800 4100 2098 4114
rect 1900 3708 2098 4100
rect 1900 3492 2096 3708
rect 1900 3400 2098 3492
rect 1945 2955 2054 3400
rect -672 2896 -480 2904
rect -1581 1325 -1575 1476
rect -1424 1325 -1418 1476
rect -1581 1313 -1418 1325
rect -2528 910 -2522 1090
rect -2342 910 -2336 1090
rect -2528 898 -2336 910
rect -1056 868 -992 2632
rect -672 2596 -480 2704
rect 1028 2896 1220 2904
rect 1945 2840 2054 2846
rect 1028 2504 1220 2704
rect -928 1490 -736 2396
rect -928 1310 -922 1490
rect -742 1310 -736 1490
rect -928 1298 -736 1310
rect 644 868 708 2132
rect 772 1490 964 2396
rect 772 1310 778 1490
rect 958 1310 964 1490
rect 1219 1399 1319 1405
rect 772 1298 964 1310
rect 1043 1393 1219 1399
rect 1043 1305 1055 1393
rect 1143 1305 1219 1393
rect 1043 1299 1219 1305
rect 1219 1293 1319 1299
<< via1 >>
rect -2481 6075 -2318 6081
rect -2481 5924 -2475 6075
rect -2475 5924 -2324 6075
rect -2324 5924 -2318 6075
rect -2481 5918 -2318 5924
rect -1581 5918 -1418 6081
rect -2272 4804 -2080 4996
rect -2656 2868 -2592 2932
rect 1004 4804 1196 4996
rect 1914 4114 2085 4285
rect -672 2704 -480 2896
rect 1028 2704 1220 2896
rect 1945 2846 2054 2955
rect 1219 1299 1319 1399
<< metal2 >>
rect -2487 5918 -2481 6081
rect -2318 5918 -1581 6081
rect -1418 5918 -1412 6081
rect 990 4996 1227 5012
rect -2278 4804 -2272 4996
rect -2080 4804 1004 4996
rect 1196 4804 1227 4996
rect 990 4791 1227 4804
rect 1908 4284 1914 4285
rect 1906 4114 1914 4284
rect 2085 4284 2091 4285
rect 2085 4114 2092 4284
rect 1906 4098 2092 4114
rect 1910 3868 2092 4098
rect 1908 3851 2334 3868
rect 1908 3717 2177 3851
rect 2311 3717 2334 3851
rect 1908 3702 2334 3717
rect -2678 2932 1945 2955
rect -2678 2868 -2656 2932
rect -2592 2896 1945 2932
rect -2592 2868 -672 2896
rect -2678 2846 -672 2868
rect -678 2704 -672 2846
rect -480 2846 1028 2896
rect -480 2704 -474 2846
rect 1022 2704 1028 2846
rect 1220 2846 1945 2896
rect 2054 2846 2060 2955
rect 1220 2704 1226 2846
rect 1386 1399 1476 1403
rect 1213 1299 1219 1399
rect 1319 1394 1481 1399
rect 1319 1304 1386 1394
rect 1476 1304 1481 1394
rect 1319 1299 1481 1304
rect 1386 1295 1476 1299
<< via2 >>
rect 2177 3717 2311 3851
rect 1386 1304 1476 1394
<< metal3 >>
rect -8700 6300 1800 6400
rect 1700 4800 1800 6300
rect -8700 4700 1800 4800
rect 1700 3500 1800 4700
rect 2160 3856 2332 3870
rect 2160 3712 2172 3856
rect 2316 3712 2332 3856
rect 2160 3700 2332 3712
rect -8700 3400 1800 3500
rect 1700 2062 1800 3400
rect 1699 2000 1800 2062
rect -8700 1900 1800 2000
rect 1699 1399 1799 1900
rect 1381 1394 1799 1399
rect 1381 1304 1386 1394
rect 1476 1304 1799 1394
rect 1381 1299 1799 1304
<< via3 >>
rect 2172 3851 2316 3856
rect 2172 3717 2177 3851
rect 2177 3717 2311 3851
rect 2311 3717 2316 3851
rect 2172 3712 2316 3717
<< metal4 >>
rect -8700 6300 1800 6400
rect 1700 4800 1800 6300
rect -8700 4700 1800 4800
rect 1700 3851 1800 4700
rect 2171 3856 2317 3857
rect 2171 3851 2172 3856
rect 1700 3717 2172 3851
rect 1700 3671 1800 3717
rect 2171 3712 2172 3717
rect 2316 3712 2317 3856
rect 2171 3711 2317 3712
rect -8700 3400 1800 3500
rect 1700 2000 1800 3400
rect -8700 1900 1800 2000
use JNWTR_CAPX1  JNWTR_CAPX1_0 ../JNW_TR_SKY130A
array 0 7 1350 0 3 1350
timestamp 1735426800
transform 1 0 -8700 0 1 1900
box 0 0 1080 1080
use JNWATR_PCH_2C5F0  x1 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 -1216 0 1 2028
box -184 -128 1208 928
use JNWATR_NCH_2C5F0  x2 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 -2816 0 1 2028
box -184 -128 1208 928
use JNWTR_RPPO16  x3 ../JNW_TR_SKY130A
timestamp 1735575823
transform 1 0 -2900 0 1 3000
box 0 0 4472 3440
use JNWATR_PCH_2C5F0  x5
timestamp 1734044400
transform 1 0 484 0 1 2028
box -184 -128 1208 928
<< labels >>
flabel locali -700 1200 778 1600 0 FreeSans 1600 0 0 0 VDD_1V8
port 1 nsew
flabel locali -3500 6600 2100 7000 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal1 644 868 708 2132 0 FreeSans 800 90 0 0 RESET_N_1V8
port 4 nsew
flabel metal1 -1056 868 -992 2328 0 FreeSans 800 90 0 0 PWRUP_B_1V8
port 5 nsew
flabel metal1 1000 5300 2100 5500 0 FreeSans 1600 0 0 0 VO_1V8
port 6 nsew
flabel metal1 1900 3400 1910 4114 0 FreeSans 1600 0 0 0 IPTN
port 3 nsew
<< end >>
