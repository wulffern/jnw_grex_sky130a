magic
tech sky130A
magscale 1 2
timestamp 1735576154
<< locali >>
rect -200 -2200 6600 -2000
rect -200 -8000 0 -2200
rect 200 -2496 6198 -2400
rect 200 -2676 4276 -2496
rect 4456 -2676 6198 -2496
rect 200 -2800 6198 -2676
rect 3886 -3257 4078 -2800
rect 4910 -3257 5102 -2800
rect 2165 -3999 2357 -3757
rect 3189 -3999 3381 -3767
rect 2165 -4005 3381 -3999
rect 2165 -4185 2555 -4005
rect 2735 -4185 3381 -4005
rect 2165 -4387 3381 -4185
rect 6400 -4387 6600 -2200
rect 1846 -4499 6600 -4387
rect 346 -8000 538 -7646
rect 1370 -8000 1562 -7598
rect 1846 -8000 1958 -7651
rect 6174 -8000 6286 -7683
rect 6400 -8000 6600 -4499
rect -200 -8122 6600 -8000
rect -200 -8302 736 -8122
rect 916 -8302 6600 -8122
rect -200 -8400 6600 -8302
<< viali >>
rect 4276 -2676 4456 -2496
rect 2555 -4185 2735 -4005
rect 2230 -4821 2410 -4641
rect 5679 -4838 5859 -4658
rect 736 -8302 916 -8122
<< metal1 >>
rect 1786 -2800 1978 -2794
rect 602 -3524 666 -3518
rect 1064 -3524 1128 -3518
rect 602 -4708 666 -3588
rect 986 -3588 1064 -3543
rect 1128 -3588 1324 -3543
rect 986 -3735 1324 -3588
rect 1516 -3735 1522 -3543
rect 1786 -3885 1978 -2992
rect 2421 -2920 2485 -2914
rect 2421 -3740 2485 -2984
rect 4142 -2917 4206 -2395
rect 2799 -3174 3009 -3168
rect 4142 -3234 4206 -2981
rect 4270 -2496 4462 -2484
rect 4270 -2676 4276 -2496
rect 4456 -2676 4462 -2496
rect 2799 -3390 3009 -3384
rect 980 -4077 986 -3885
rect 1178 -4077 1184 -3885
rect 1786 -4083 1978 -4077
rect 2549 -4005 2741 -3575
rect 4270 -3616 4462 -2676
rect 2549 -4185 2555 -4005
rect 2735 -4185 2741 -4005
rect 2549 -4197 2741 -4185
rect 4526 -4090 4718 -3583
rect 732 -4294 924 -4288
rect 732 -4492 924 -4486
rect 1308 -4294 1534 -4284
rect 4526 -4288 4718 -4282
rect 5673 -4090 5865 -4084
rect 1308 -4486 1320 -4294
rect 1512 -4486 1534 -4294
rect 1308 -4496 1534 -4486
rect 602 -5190 666 -4772
rect 1070 -4708 1134 -4702
rect 1070 -4778 1134 -4772
rect 736 -4952 928 -4946
rect 736 -5150 928 -5144
rect 1070 -5518 1134 -5512
rect 1070 -5588 1134 -5582
rect 602 -7126 666 -6008
rect 602 -7262 666 -7190
rect 730 -8122 922 -5820
rect 1320 -6338 1512 -4496
rect 2218 -4504 2224 -4312
rect 2416 -4504 2422 -4312
rect 2224 -4641 2416 -4504
rect 2224 -4821 2230 -4641
rect 2410 -4821 2416 -4641
rect 2224 -4833 2416 -4821
rect 5673 -4658 5865 -4282
rect 5673 -4838 5679 -4658
rect 5859 -4838 5865 -4658
rect 5673 -4850 5865 -4838
rect 1320 -6536 1512 -6530
rect 1058 -7126 1122 -7120
rect 1058 -7196 1122 -7190
rect 730 -8302 736 -8122
rect 916 -8302 922 -8122
rect 730 -8314 922 -8302
<< via1 >>
rect 1786 -2992 1978 -2800
rect 730 -3380 922 -3188
rect 602 -3588 666 -3524
rect 1064 -3588 1128 -3524
rect 1324 -3735 1516 -3543
rect 2421 -2984 2485 -2920
rect 4142 -2981 4206 -2917
rect 2799 -3384 3009 -3174
rect 986 -4077 1178 -3885
rect 1786 -4077 1978 -3885
rect 4526 -4282 4718 -4090
rect 732 -4486 924 -4294
rect 5673 -4282 5865 -4090
rect 1320 -4486 1512 -4294
rect 602 -4772 666 -4708
rect 1070 -4772 1134 -4708
rect 736 -5144 928 -4952
rect 602 -5582 666 -5518
rect 1070 -5582 1134 -5518
rect 602 -7190 666 -7126
rect 2224 -4504 2416 -4312
rect 986 -6530 1178 -6338
rect 1320 -6530 1512 -6338
rect 1058 -7190 1122 -7126
<< metal2 >>
rect 1766 -2800 1992 -2788
rect 1766 -2992 1786 -2800
rect 1978 -2992 1992 -2800
rect 4137 -2917 4214 -2908
rect 2291 -2920 4142 -2917
rect 2291 -2981 2421 -2920
rect 2415 -2984 2421 -2981
rect 2485 -2981 4142 -2920
rect 4206 -2981 4214 -2917
rect 2485 -2984 2491 -2981
rect 1766 -3010 1992 -2992
rect 4137 -2995 4214 -2981
rect 261 -3188 2799 -3174
rect 261 -3380 280 -3188
rect 472 -3380 730 -3188
rect 922 -3380 2799 -3188
rect 261 -3384 2799 -3380
rect 3009 -3384 3015 -3174
rect 578 -3524 678 -3508
rect 1060 -3524 1160 -3508
rect 578 -3588 602 -3524
rect 666 -3588 1064 -3524
rect 1128 -3588 1160 -3524
rect 578 -3602 678 -3588
rect 1060 -3602 1160 -3588
rect 1324 -3543 1516 -3537
rect 1516 -3735 2408 -3543
rect 1324 -3741 1516 -3735
rect 986 -3885 1178 -3879
rect 1178 -4077 1786 -3885
rect 1978 -4077 1984 -3885
rect 986 -4083 1178 -4077
rect 2216 -4268 2408 -3735
rect 1308 -4294 1534 -4284
rect 726 -4486 732 -4294
rect 924 -4486 1320 -4294
rect 1512 -4486 1534 -4294
rect 1308 -4496 1534 -4486
rect 2216 -4312 2416 -4268
rect 4520 -4282 4526 -4090
rect 4718 -4282 5673 -4090
rect 5865 -4282 5871 -4090
rect 2216 -4504 2224 -4312
rect 2216 -4506 2416 -4504
rect 2224 -4510 2416 -4506
rect 580 -4708 680 -4692
rect 1056 -4708 1156 -4686
rect 580 -4772 602 -4708
rect 666 -4772 1070 -4708
rect 1134 -4772 1156 -4708
rect 580 -4786 680 -4772
rect 1056 -4780 1156 -4772
rect 280 -4957 736 -4952
rect 276 -5139 285 -4957
rect 467 -5139 736 -4957
rect 280 -5144 736 -5139
rect 928 -5144 934 -4952
rect 582 -5518 682 -5504
rect 1056 -5518 1156 -5498
rect 295 -5582 304 -5518
rect 368 -5582 602 -5518
rect 666 -5582 1070 -5518
rect 1134 -5582 1156 -5518
rect 582 -5598 682 -5582
rect 1056 -5592 1156 -5582
rect 974 -6338 1190 -6324
rect 974 -6530 986 -6338
rect 1178 -6530 1320 -6338
rect 1512 -6530 1518 -6338
rect 974 -6541 1190 -6530
rect 590 -7126 682 -7116
rect 590 -7190 602 -7126
rect 666 -7190 1058 -7126
rect 1122 -7190 1128 -7126
rect 590 -7196 682 -7190
<< via2 >>
rect 1786 -2992 1978 -2800
rect 280 -3380 472 -3188
rect 285 -5139 467 -4957
rect 304 -5582 368 -5518
<< metal3 >>
rect 1786 -2795 1978 -1854
rect 1781 -2800 1983 -2795
rect 1781 -2992 1786 -2800
rect 1978 -2992 1983 -2800
rect 1781 -2997 1983 -2992
rect 275 -3188 477 -3183
rect 275 -3380 280 -3188
rect 472 -3380 477 -3188
rect 275 -3385 477 -3380
rect 280 -4957 472 -3385
rect 280 -5139 285 -4957
rect 467 -5139 472 -4957
rect 280 -5518 472 -5139
rect 280 -5582 304 -5518
rect 368 -5582 472 -5518
rect 280 -5798 472 -5582
use JNWATR_NCH_2C5F0  JNWATR_NCH_2C5F0_0 ../JNW_ATR_SKY130A
array 0 0 1024 0 5 800
timestamp 1734044400
transform 1 0 442 0 1 -7798
box -184 -128 1208 928
use JNWATR_NCH_2C5F0  x1
timestamp 1734044400
transform 1 0 2261 0 1 -3920
box -184 -128 1208 928
use JNWTR_RPPO16  x3 ../JNW_TR_SKY130A
timestamp 1735575823
transform 1 0 1830 0 1 -7811
box 0 0 4472 3440
use JNWATR_PCH_2C1F2  x4 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 3982 0 1 -3905
box -184 -128 1208 928
<< labels >>
flabel metal3 280 -4957 472 -3380 0 FreeSans 640 90 0 0 VBN2
flabel metal1 4142 -3405 4206 -2395 0 FreeSans 800 90 0 0 PWRUP_N_1V8
port 5 nsew
flabel locali 200 -2800 4276 -2400 0 FreeSans 1600 0 0 0 VDD_1V8
port 7 nsew
flabel locali 916 -8400 6600 -8000 0 FreeSans 1600 0 0 0 VSS
port 8 nsew
flabel metal3 1786 -2800 1978 -1854 0 FreeSans 1600 90 0 0 IPTN
<< end >>
