*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/JNWGREX_TI_lpe.spi
#else
.include ../../../work/xsch/JNWGREX_TI.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
*.option TNOM=27 GMIN=1e-15 reltol=1e-3
.option reltol=1e-4
*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  0 dc {AVDD}
VPWR PWRUP_N_1V8 0 dc 0


VO IPTN 0 dc 0.9

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all

B5 temp 0 v=temper

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 100n 10u 0


dc TEMP -40 100 5

print v(temp-sweep)


let vbn2_d1 = deriv(v(xdut.vbn2))/deriv(v(temp))
let vbn2_d2 = deriv(vbn2_d1)/deriv(v(temp))

write
quit


.endc

.end
