magic
tech sky130A
magscale 1 2
timestamp 1735576154
<< locali >>
rect -400 6300 14800 6500
rect -400 5800 -200 6300
rect 14298 3763 14474 3769
rect 14298 3599 14304 3763
rect 14468 3599 14474 3763
rect 14298 2730 14474 3599
rect 14290 2675 14474 2730
rect 12727 2370 12979 2430
rect 12919 2030 12979 2370
rect 14290 2155 14461 2675
rect 12919 1970 13270 2030
rect 13821 1876 14107 1926
rect 12730 1263 12790 1559
rect 13821 1553 13871 1876
rect 13710 1503 13871 1553
rect 12887 1230 12947 1329
rect 12887 1170 13091 1230
rect 13813 1089 14039 1141
rect 12615 910 12984 957
rect 12615 897 13090 910
rect 13813 902 13865 1089
rect 12924 850 13090 897
rect 13709 850 13865 902
rect 12877 606 12977 666
rect 12917 590 12977 606
rect 12917 530 13418 590
rect 13787 440 14109 500
rect 12589 270 12967 325
rect 13787 270 13847 440
rect 12589 265 13090 270
rect 12907 210 13090 265
rect 13449 210 13847 270
rect 12309 -200 12491 91
rect -400 -359 12792 -200
rect 14600 -200 14800 6300
rect 12956 -359 14800 -200
rect -400 -400 14800 -359
<< viali >>
rect 2597 5200 2997 5600
rect 9665 5000 10065 5400
rect 14304 3599 14468 3763
rect 13400 2626 13449 2675
rect 12756 2564 12804 2612
rect 13332 1958 13392 2018
rect 12730 1203 12790 1263
rect 12887 1329 12947 1389
rect 12555 897 12615 957
rect 13930 700 14030 800
rect 12817 606 12877 666
rect 12529 265 12589 325
rect 13936 106 14024 194
rect 12792 -359 12956 -195
<< metal1 >>
rect 12692 6182 12756 6188
rect 8844 6070 8908 6076
rect 3942 6022 4006 6028
rect 2597 5817 2997 5823
rect 2580 5200 2597 5612
rect 2997 5200 3049 5612
rect 2580 5179 3049 5200
rect 3942 5117 4006 5958
rect 12424 6006 12430 6070
rect 12494 6006 12500 6070
rect 8844 5668 8908 6006
rect 10544 5862 10608 5868
rect 9665 5852 10065 5858
rect 10544 5668 10608 5798
rect 12430 5746 12494 6006
rect 12331 5682 12494 5746
rect 12546 5862 12610 5868
rect 9665 5406 10065 5452
rect 12107 5646 12276 5652
rect 9653 5400 10077 5406
rect 9653 5000 9665 5400
rect 10065 5000 10077 5400
rect 9653 4994 10077 5000
rect 12107 3775 12276 5477
rect 12107 3769 12283 3775
rect 12107 3587 12283 3593
rect 12107 3558 12276 3587
rect 12127 2618 12187 2624
rect 11713 1263 11997 1292
rect 11713 1232 11776 1263
rect 11836 1232 11997 1263
rect 11776 1197 11836 1203
rect 12127 666 12187 2558
rect 12331 1406 12395 5682
rect 12546 5570 12610 5798
rect 12438 5506 12610 5570
rect 12307 1389 12407 1406
rect 12307 1329 12329 1389
rect 12389 1329 12407 1389
rect 12307 1320 12407 1329
rect 12127 600 12187 606
rect 12438 340 12502 5506
rect 12692 5384 12756 6118
rect 12552 5320 12756 5384
rect 12552 969 12616 5320
rect 14298 3769 14474 3775
rect 14298 3587 14474 3593
rect 14200 2681 14500 2700
rect 13388 2675 14500 2681
rect 13388 2626 13400 2675
rect 13449 2626 14500 2675
rect 12750 2618 12810 2624
rect 13388 2620 14500 2626
rect 14200 2600 14500 2620
rect 12750 2552 12810 2558
rect 13320 2018 14012 2024
rect 13320 1958 13332 2018
rect 13392 2000 14012 2018
rect 13392 1958 14500 2000
rect 13320 1952 14500 1958
rect 13926 1900 14500 1952
rect 12875 1389 12893 1395
rect 12875 1329 12887 1389
rect 12875 1323 12893 1329
rect 12953 1323 12959 1395
rect 12711 1269 12811 1275
rect 12711 1197 12724 1269
rect 12796 1197 12811 1269
rect 12711 1190 12811 1197
rect 12549 957 12621 969
rect 12549 897 12555 957
rect 12615 897 12621 957
rect 12549 885 12621 897
rect 12552 809 12616 885
rect 13918 800 14042 806
rect 13918 700 13930 800
rect 14030 700 14500 800
rect 13918 694 14042 700
rect 12811 672 12883 678
rect 12805 600 12811 672
rect 12871 666 12883 672
rect 12877 606 12883 666
rect 12871 600 12883 606
rect 12811 594 12883 600
rect 12438 325 12595 340
rect 12436 265 12529 325
rect 12589 265 12595 325
rect 12438 239 12595 265
rect 12438 202 12502 239
rect 13924 194 14500 200
rect 13924 106 13936 194
rect 14024 106 14500 194
rect 13924 100 14500 106
rect 12780 -195 13030 -189
rect 12780 -359 12792 -195
rect 12956 -359 13030 -195
rect 12780 -365 13030 -359
rect 13206 -365 13212 -189
<< via1 >>
rect 12692 6118 12756 6182
rect 3942 5958 4006 6022
rect 2597 5600 2997 5817
rect 2597 5417 2997 5600
rect 8844 6006 8908 6070
rect 12430 6006 12494 6070
rect 9665 5452 10065 5852
rect 10544 5798 10608 5862
rect 12546 5798 12610 5862
rect 12107 5477 12276 5646
rect 12107 3593 12283 3769
rect 12127 2558 12187 2618
rect 11776 1203 11836 1263
rect 12329 1329 12389 1389
rect 12127 606 12187 666
rect 14298 3763 14474 3769
rect 14298 3599 14304 3763
rect 14304 3599 14468 3763
rect 14468 3599 14474 3763
rect 14298 3593 14474 3599
rect 12750 2612 12810 2618
rect 12750 2564 12756 2612
rect 12756 2564 12804 2612
rect 12804 2564 12810 2612
rect 12750 2558 12810 2564
rect 12893 1389 12953 1395
rect 12893 1329 12947 1389
rect 12947 1329 12953 1389
rect 12893 1323 12953 1329
rect 12724 1263 12796 1269
rect 12724 1203 12730 1263
rect 12730 1203 12790 1263
rect 12790 1203 12796 1263
rect 12724 1197 12796 1203
rect 12811 666 12871 672
rect 12811 606 12817 666
rect 12817 606 12871 666
rect 12811 600 12871 606
rect 13030 -365 13206 -189
<< metal2 >>
rect 1603 6150 1612 6259
rect 1721 6254 6270 6259
rect 1721 6155 6166 6254
rect 6265 6155 6274 6254
rect 1721 6150 6270 6155
rect 8649 6118 12692 6182
rect 12756 6118 12762 6182
rect 8649 6022 8713 6118
rect 12430 6070 12494 6076
rect 3936 5958 3942 6022
rect 4006 5958 8713 6022
rect 8838 6006 8844 6070
rect 8908 6006 12430 6070
rect 12430 6000 12494 6006
rect 1 5852 10071 5858
rect 1 5817 9665 5852
rect 1 5446 2597 5817
rect 2580 5417 2597 5446
rect 2997 5452 9665 5817
rect 10065 5646 10071 5852
rect 10538 5798 10544 5862
rect 10608 5798 12546 5862
rect 12610 5798 12616 5862
rect 10065 5477 12107 5646
rect 12276 5477 12282 5646
rect 10065 5452 10071 5477
rect 2997 5446 10071 5452
rect 2997 5417 3049 5446
rect 2580 5179 3049 5417
rect 6188 5088 6297 5097
rect 6188 3754 6297 4979
rect 13575 3769 13741 3773
rect 6188 3645 8156 3754
rect 12101 3593 12107 3769
rect 12283 3764 14298 3769
rect 12283 3598 13575 3764
rect 13741 3598 14298 3764
rect 12283 3593 14298 3598
rect 14474 3593 14480 3769
rect 13575 3589 13741 3593
rect 12121 2558 12127 2618
rect 12187 2558 12750 2618
rect 12810 2558 12816 2618
rect 12893 1395 12953 1401
rect 12323 1329 12329 1389
rect 12389 1329 12893 1389
rect 12893 1317 12953 1323
rect 12711 1269 12811 1275
rect 12711 1263 12724 1269
rect 11770 1203 11776 1263
rect 11836 1203 12724 1263
rect 12711 1197 12724 1203
rect 12796 1197 12811 1269
rect 12711 1190 12811 1197
rect 12811 672 12871 678
rect 12121 606 12127 666
rect 12187 606 12811 666
rect 12811 594 12871 600
rect 13030 -104 13206 -99
rect 13026 -189 13035 -104
rect 13201 -189 13210 -104
rect 13026 -270 13030 -189
rect 13206 -270 13210 -189
rect 13030 -371 13206 -365
<< via2 >>
rect 1612 6150 1721 6259
rect 6166 6155 6265 6254
rect 6188 4979 6297 5088
rect 13575 3598 13741 3764
rect 13035 -189 13201 -104
rect 13035 -270 13201 -189
<< metal3 >>
rect 1607 6259 1726 6264
rect 1607 6150 1612 6259
rect 1721 6150 1726 6259
rect 1607 6145 1726 6150
rect 6154 6254 6306 6266
rect 6154 6155 6166 6254
rect 6265 6155 6306 6254
rect 1612 5621 1721 6145
rect 6154 6136 6306 6155
rect 6188 5093 6297 6136
rect 6183 5088 6302 5093
rect 6183 4979 6188 5088
rect 6297 4979 6302 5088
rect 6183 4974 6302 4979
rect 13570 3764 13746 3769
rect 6156 3640 6161 3759
rect 6270 3640 6275 3759
rect 13570 3598 13575 3764
rect 13741 3598 13746 3764
rect 13570 2864 13746 3598
rect 13030 -104 13206 1341
rect 13574 251 13743 2730
rect 13030 -270 13035 -104
rect 13201 -270 13206 -104
rect 13030 -275 13206 -270
use JNWTR_TAPCELLB_CV  JNWTR_TAPCELLB_CV_0 ~/data/2023/aicex/ip/jnw_grex_sky130a/design/JNW_TR_SKY130A
timestamp 1735485359
transform 1 0 12400 0 1 2720
box -150 -120 2130 440
use JNWGREX_TI  XA_TI1
timestamp 1735576154
transform 1 0 -200 0 1 8000
box -200 -8400 6600 -1854
use JNWGREX_ITD  XB_ITD1
timestamp 1735576154
transform 1 0 9900 0 -1 6600
box -8700 868 2100 7030
use JNWTR_IVX1_CV  xc1 ~/data/2023/aicex/ip/jnw_grex_sky130a/design/JNW_GREX_SKY130A/../JNW_TR_SKY130A
timestamp 1735576154
transform 1 0 12400 0 1 0
box -150 -120 2130 440
use JNWTR_IVX1_CV  xc2
timestamp 1735576154
transform 1 0 12400 0 1 320
box -150 -120 2130 440
use JNWTR_IVX1_CV  xc3
timestamp 1735576154
transform 1 0 12400 0 1 640
box -150 -120 2130 440
use JNWTR_IVX1_CV  xc4
timestamp 1735576154
transform 1 0 12400 0 1 960
box -150 -120 2130 440
use JNWTR_IVX2_CV  xc5 ~/data/2023/aicex/ip/jnw_grex_sky130a/design/JNW_GREX_SKY130A/../JNW_TR_SKY130A
timestamp 1735576154
transform 1 0 12400 0 1 1280
box -150 -120 2130 600
use JNWTR_IVX2_CV  xc6
timestamp 1735576154
transform 1 0 12400 0 1 1760
box -150 -120 2130 600
use JNWTR_NRX1_CV  xc7 ~/data/2023/aicex/ip/jnw_grex_sky130a/design/JNW_GREX_SKY130A/../JNW_TR_SKY130A
timestamp 1735576154
transform 1 0 12400 0 1 2240
box -150 -120 2130 600
<< labels >>
flabel space 13030 210 13847 270 0 FreeSans 480 0 0 0 RESET_N_1V8
flabel space 13030 530 13660 590 0 FreeSans 480 0 0 0 RESET_B_1V8
flabel space 13030 850 13660 910 0 FreeSans 480 0 0 0 PWRUP_N_1V8
flabel space 13030 1170 13660 1230 0 FreeSans 480 0 0 0 PWRUP_B_1V8
flabel space 13030 1490 13660 1550 0 FreeSans 480 0 0 0 VO_N_1V8
flabel space 13270 2610 13660 2670 0 FreeSans 480 0 0 0 PULSE_1V8
port 3 nsew
flabel metal1 14200 2600 14500 2700 0 FreeSans 640 0 0 0 PULSE_1V8
port 6 nsew
flabel metal1 14200 1900 14500 2000 0 FreeSans 640 0 0 0 DO_1V8
port 7 nsew
flabel metal1 14200 700 14500 800 0 FreeSans 640 0 0 0 PWRUP_1V8
port 8 nsew
flabel metal1 14200 100 14500 200 0 FreeSans 640 0 0 0 RESET_1V8
port 9 nsew
flabel metal2 1 5446 413 5858 0 FreeSans 1600 90 0 0 VDD_1V8
port 4 nsew
flabel locali -400 -400 12792 -200 0 FreeSans 1600 0 0 0 VSS
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 14380 6400
<< end >>
